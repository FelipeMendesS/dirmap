----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    10:51:17 11/02/2016 
-- Design Name: 
-- Module Name:    aux_control_cell - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity aux_control_cell is
    Port ( Ri : in  STD_LOGIC;
           Ai : in  STD_LOGIC;
           Ro : out  STD_LOGIC;
           Ao : out  STD_LOGIC);
end aux_control_cell;

architecture Behavioral of aux_control_cell is

begin


end Behavioral;

